//rising edge detector

module rising_edge();
	
	
endmodule

